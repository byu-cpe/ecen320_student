/***************************************************************************
* 
* Filename: logic_functions.sv
*
* Author: <Your Name>
* Description: <Provide a description of what this HDL file does>
*
****************************************************************************/

module logic_functions (
        input logic     A,
        input logic     B,
        input logic     C,
        output logic    O1,
        output logic    O2
    );

// O1 = AC+A'B

// O2 = (A+C')(BC)

endmodule